`timescale 1ns/1ns


module datapath_tb;
    reg [31:0]intTr;
    wire TR_ZF;


datapath DUV(intTr,TR_ZF);

initial 
begin
    $dumpfile("datapath_tb.vcd");
    $dumpvars(0,datapath_tb);

    //ADD         
    #100;intTr=32'b00000000111010100100000000100000;//8
    #100;intTr=32'b00000010010010100100100000100000;//9
    
    //AND
    #100;intTr=32'b00000000010010110101000000100100;//10
    #100;intTr=32'b00000011111110100101100000100100;//11

    //SUB
    #100;intTr=32'b00000011110101000110000000100010;//12
    #100;intTr=32'b00000000011011110110100000100010;//13

    //OR
    #100;intTr=32'b00000010001001110111000000100101;//14
    #100;intTr=32'b00000010101010110111100000100101;//15

    //SLT
    #100;intTr=32'b00000010000101001000000000100101;//16
    #100;intTr=32'b00000011101000101000100000100101;//17
    $stop;
end

endmodule